// module flipflop(
//     clk,
//     rst_n,
//     CurrentState,
//     NextState,
// );
// input clk; 
// input rst_n;
// input CurrentState;
// output NextState;


// always @(posedge clk or negedge rst_n)
// begin
//     if(!rst_n)
//     CurrentState <= green_h;
//     else 
//     CurrentState <= NextState;
// end

// endmodule